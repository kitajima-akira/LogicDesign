// decoder_7seg_table.sv - 7セグメントLEDデコーダ (テーブル方式)

//! 7セグメントLEDデコーダ
//
//        --y[6]--
//       /        /
//     y[1]      y[5]
//      /        /
//      /--y[0]--/
//      /        /
//    y[2]     y[4]
//     /        /
//      --y[3]--
module decoder_7seg_table(
    input logic[3:0] d,  //! 入力値
    output logic[6:0] y  //! 対応する7セグメントLEDの点灯パターン
  );

  always_comb
  begin
    case(d)
      'b0000:
        y = 'b1111110; // 0
      'b0001:
        y = 'b0110000; // 1
      'b0010:
        y = 'b1101101; // 2
      'b0011:
        y = 'b1111001; // 3
      'b0100:
        y = 'b0110011; // 4
      'b0101:
        y = 'b1011011; // 5
      'b0110:
        y = 'b1011111; // 6
      'b0111:
        y = 'b1110000; // 7
      'b1000:
        y = 'b1111111; // 8
      'b1001:
        y = 'b1111011; // 9
      'b1010:
        y = 'b1110111; // A
      'b1011:
        y = 'b0011111; // b
      'b1100:
        y = 'b1001110; // C
      'b1101:
        y = 'b0111101; // d
      'b1110:
        y = 'b1001111; // E
      'b1111:
        y = 'b1000111; // F
      default:
        y = 'b1111111; // その他
    endcase
  end
endmodule
