// full_adder_tb.sv - 全加算器のテストベンチ

// 全加算器のテストベンチ
module full_adder_tb;
  // 入力用信号
  logic a;
  logic b;
  logic ci;

  // 出力用信号
  logic s;
  logic co;

  // テスト対象回路 UUT (the Unit Under Test)
  full_adder uut(.*);

  // 波形生成
  initial
  begin
    // ヘッダ表示
    $display("a b ci:co s");
    $display("- - - + - -");

    // テストパターンの生成 (全組み合わせ)
    for (int i = 0; i < 8; i++)
    begin
      a = i[2];
      b = i[1];
      ci = i[0];

      #10
       $display("%b %b %b : %b %b", a, b, ci, co, s);
    end

    // シミュレーション終了
    $finish;
  end
endmodule
